module calculadora (
    input logic [3] cmd,
    input logic clock,
    input logic reset,
    
    output logic [1] status,
    output logic [3] data,
    output logic [3] position
);
    
endmodule