module calculadora (
    input logic [3] cmd,
    input logic clock,
    input logic reset,
    
    output logic [2] status,
    output logic [4] data,
    output logic [4] position
);
    
endmodule